`define x1 0
`define x2 0
`define x3 1
`define x4 1
`define x5 2
`define x6 2
`define x7 2
`define x8 2
`define x9 2
`define x10 2
`define x11 2
`define x12 2
`define x13 2
`define x14 2
`define x15 3
`define x16 3
`define x17 4
`define x18 4
`define x19 5
`define x20 5
`define x21 6
`define x22 6
`define x23 6

`define y1 3
`define y2 4
`define y3 1
`define y4 2
`define y5 0
`define y6 1
`define y7 2
`define y8 3
`define y9 4
`define y10 5
`define y11 6
`define y12 7
`define y13 8
`define y14 9
`define y15 6
`define y16 9
`define y17 5
`define y18 9
`define y19 5
`define y20 9
`define y21 6
`define y22 7
`define y23 8
