`define x1 0
`define x2 0
`define x3 0
`define x4 1
`define x5 1
`define x6 1
`define x7 1
`define x8 1
`define x9 2
`define x10 2
`define x11 2
`define x12 2
`define x13 3
`define x14 3
`define x15 3
`define x16 4
`define x17 4
`define x18 4
`define x19 5
`define x20 5
`define x21 5
`define x22 5
`define x23 5
`define x24 5
`define x25 5
`define x26 5
`define x27 5
`define x28 5
`define x29 5
`define x30 5
`define x31 5
`define x32 5
`define x33 5
`define x34 5
`define x35 5
`define x36 6
`define x37 6
`define x38 6
`define x39 6
`define x40 7
`define x41 7
`define x42 8
`define x43 8
`define x44 8
`define x45 8
`define x46 9
`define x47 9
`define x48 9
`define x49 10
`define x50 10
`define x51 10
`define x52 11
`define x53 11
`define x54 11
`define x55 12
`define x56 12
`define x57 12
`define x58 12
`define x59 13
`define x60 13
`define x61 14
`define x62 14
`define x63 14
`define x64 14
`define x65 14


`define y1 5
`define y2 6
`define y3 7
`define y4 4
`define y5 5
`define y6 6
`define y7 7
`define y8 8
`define y9 3
`define y10 4
`define y11 5
`define y12 9
`define y13 2
`define y14 3
`define y15 4
`define y16 1
`define y17 2
`define y18 3
`define y19 0
`define y20 1
`define y21 2
`define y22 3
`define y23 4
`define y24 5
`define y25 6
`define y26 7
`define y27 8
`define y28 9
`define y29 10
`define y30 11
`define y31 12
`define y32 13
`define y33 14
`define y34 15
`define y35 16
`define y36 11
`define y37 12
`define y38 15
`define y39 16
`define y40 10
`define y41 17
`define y42 10
`define y43 12
`define y44 13
`define y45 17
`define y46 9
`define y47 15
`define y48 17
`define y49 9
`define y50 15
`define y51 17
`define y52 9
`define y53 15
`define y54 17
`define y55 10
`define y56 12
`define y57 13
`define y58 17
`define y59 10
`define y60 16
`define y61 11
`define y62 12
`define y63 13
`define y64 14
`define y65 15
